module nnoc ();
endmodule
