module cnn ();

endmodule
